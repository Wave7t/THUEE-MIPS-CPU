`timescale 1ns/1ps

`include "defs.v"


module ID_stage (
    input wire clk,
    input wire reset,

    //==============================================================//
    // This stage needs not to be flushed, only hold is needed
    input wire          e_IFIDHold,
    // Write Back-Related
    input wire          e_RegWrite,
    input wire [4:0]    e_WBAddr,
    input wire [31:0]   e_WBData,

    // flow control: only j and jal instructions
    output wire         e_jump,
    output wire [31:0]  e_jumpDesti,
    // below: for Load-Use hanzard detection
    output wire         e_UseData1,
    output wire         e_UseData2,
    output wire [4:0]   e_rs,
    output wire [4:0]   e_rt,
`ifdef OPT_3
    input wire          e_IFID_clean,
`endif

    //==============================================================//
    // pipeline inputs
    input wire [31:0] inst_i,
    input wire [31:0] pcp4_i,

    // pipeline outputs
    output wire [31:0] pcp4_o,
    output wire [31:0] regdata1_o,
    output wire [31:0] regdata2_o,
    output wire [31:0] imm32_o,
    output wire [4:0] rs_o,
    output wire [4:0] rt_o,
    output wire [4:0] rd_o,
    output wire [4:0] shamt_o,

    //==============================================================//
    // control signal pipeline outputs
    // ALU options (EX stage)

    output wire        c_AluSrc1_o,
    output wire        c_AluSrc2_o,
    output wire [4:0]  c_aluop_o,

    // flow control signals (EX stage)
    output wire [2:0]  c_BranchOption_o,
    output wire        c_jumpReg_o,

    // Write Back signals (EX, MEM and WB)
    output wire        c_WBSrc1_o,
    output wire        c_WBSrc2_o,
    output wire [1:0]  c_RegDst_o,
    output wire        c_RegWrite_o,

    // memory options (MEM stage)
    output wire [1:0]  c_MemRdOp_o,
    output wire [1:0]  c_MemWrOp_o,
    output wire        c_MemRdSign_o
    

);

    // register update
    reg [31:0] inst_reg;
    reg [31:0] pcp4_reg;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            inst_reg <= 32'b0;
            pcp4_reg <= 32'b0;
        end
`ifdef OPT_3
        else if (e_IFID_clean) begin
            inst_reg <= 32'b0;
            pcp4_reg <= 32'b0;
        end
`endif
        else if (~e_IFIDHold) begin
            inst_reg <= inst_i;
            pcp4_reg <= pcp4_i;
        end
    end

    // components of instruction
    wire [5:0]  opcode   = inst_reg[31:26];
    wire [4:0]  rs       = inst_reg[25:21];
    wire [4:0]  rt       = inst_reg[20:16];
    wire [4:0]  rd       = inst_reg[15:11];
    wire [4:0]  shamt    = inst_reg[10:6];
    wire [5:0]  funccode = inst_reg[5:0];
    wire [15:0] imm16    = inst_reg[16:0];


    // extrapolated immediate number
    wire [31:0] imm32;


    // control signals (generated by decoder)
    wire [1:0]  c_AluSrc1;
    wire        c_AluSrc2; 
    wire [4:0]  c_aluop;

    wire [2:0]  c_BranchOption; 
    wire        c_jumpReg;         

    wire        c_jump;         // output
    wire        c_immExtOp;     // this stage

    wire        c_WBSrc1;
    wire        c_WBSrc2;
    wire [1:0]  c_RegDst;
    wire        c_RegWrite;

    wire [1:0]  c_MemRdOp;
    wire [1:0]  c_MemWrOp;
    wire        c_MemRdSign;


    // control signal pipeline outputs
    assign c_AluSrc1_o      = c_AluSrc1[0];
    assign c_AluSrc2_o      = c_AluSrc2;
    assign c_aluop_o        = c_aluop;

    assign c_BranchOption_o = c_BranchOption;
    assign c_jumpReg_o      = c_jumpReg;

    assign c_WBSrc1_o       = c_WBSrc1;
    assign c_WBSrc2_o       = c_WBSrc2;
    assign c_RegDst_o       = c_RegDst;
    assign c_RegWrite_o     = c_RegWrite;

    assign c_MemRdOp_o      = c_MemRdOp;
    assign c_MemWrOp_o      = c_MemWrOp;
    assign c_MemRdSign_o    = c_MemRdSign;


    // instruction decoder
    mips_decoder dec (
        .opcode_i(opcode),
        .funccode_i(funccode),
        .rt0_i(rt[0]),
        .rt4_i(rt[4]),

        .c_immExtOp(c_immExtOp),
        .c_AluSrc1(c_AluSrc1),
        .c_AluSrc2(c_AluSrc2),
        .c_aluop(c_aluop),

        .c_BranchOption(c_BranchOption),
        .c_jump(c_jump),
        .c_jumpReg(c_jumpReg),

        .c_RegDst(c_RegDst),
        .c_WBSrc1(c_WBSrc1),
        .c_WBSrc2(c_WBSrc2),
        .c_RegWrite(c_RegWrite),

        .c_MemRdOp(c_MemRdOp),
        .c_MemWrOp(c_MemWrOp),
        .c_MemRdSign(c_MemRdSign),

        .use_data1(e_UseData1),
        .use_data2(e_UseData2)
    );


    // regfile IO interface
    wire [4:0] addr1_r = rs;
    wire [4:0] addr2_r = rt;
    wire [31:0] rdata1;
    wire [31:0] rdata2;


    // flow control: jump and branch can not appear simultaneously
    assign e_jump = c_jump;
    assign e_jumpDesti = {pcp4_reg[31:28],inst_reg[25:0],2'b00};
    assign e_rs = rs;
    assign e_rt = rt;
    // note UseData1 and 2 are directly connected to decoder


    // pipeline output conf
    assign pcp4_o = pcp4_reg;
    assign regdata1_o = rdata1;
    assign regdata2_o = rdata2;
    assign imm32_o = imm32;
    assign rs_o = rs;
    assign rt_o = rt;
    assign rd_o = rd;
    assign shamt_o = c_AluSrc1[1] ? 5'b10000 : shamt;


    RF1 regfile (
        .clk(clk),
        .reset(reset),
        .c_wr(e_RegWrite),
        .addr1_r(addr1_r),
        .addr2_r(addr2_r),
        .data1_o(rdata1),
        .data2_o(rdata2),
        .addr_w(e_WBAddr),
        .data_i(e_WBData)
    );

    immProc immprocessor (
        .imm16_i(imm16),
        .option(c_immExtOp),
        .imm32_o(imm32)
    );

endmodule



module immProc (
    input wire [15:0] imm16_i,
    input wire option,
    output reg [31:0] imm32_o
);
    always @(*) begin
        if (option) 
            imm32_o[31:16] <= imm16_i[15] ? 16'b11111111_11111111 : 16'b0;
        else   
            imm32_o[31:16] <= 16'b0;

        imm32_o[15:0] <= imm16_i;
    end

endmodule



// module BranchingProc (
//     input wire [31:0] data1,
//     input wire [31:0] data2,
//     input wire [2:0] branch_option,

//     output reg branch
// );
//     // 5 types of branches in total:
//     // branch on:  
//     //      Equal
//     //      Unequal
//     //      Greater than 0
//     //      Greater of Equal to 0
//     //      Less than 0
//     // And in some case, links

//     wire equal          = (data1     == data2);
//     wire is_zero        = (data1     == 32'b0);
//     wire is_negative    = (data1[31] == 1'b1);

//     always @(*) begin
//         case (branch_option) 
//             `BO_beq:    branch <= equal;
//             `BO_gez:    branch <= ~is_negative;
//             `BO_gtz:    branch <= ~(is_zero || is_negative);
//             `BO_ltz:    branch <= is_negative;
//             `BO_ueq:    branch <= ~equal;
//             `BO_lez:    branch <= is_zero || is_negative;
//             `BO_none:   branch <= 1'b0;
//             default:    branch <= 1'b0;
//         endcase
//     end
    
// endmodule



module LoadUseHanzardDetector_wo_wt (
    input wire EX_is_load,
    input wire ID_use_data1,
    input wire ID_use_data2,

    input wire [4:0] ID_raddr1,
    input wire [4:0] ID_raddr2,
    input wire [4:0] EX_waddr,

    output reg stall
);

    always @(*) begin
        if (    EX_is_load && EX_waddr != 5'b0 && 
                (
                    (ID_use_data1 && (ID_raddr1 == EX_waddr)) || 
                    (ID_use_data2 && (ID_raddr2 == EX_waddr))
                )   )
            stall <= 1'b1; 
        else 
            stall <= 1'b0;
    end
    
endmodule

